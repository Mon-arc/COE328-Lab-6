library verilog;
use verilog.vl_types.all;
entity ALU3_vlg_vec_tst is
end ALU3_vlg_vec_tst;
