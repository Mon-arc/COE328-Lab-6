library verilog;
use verilog.vl_types.all;
entity Circuit3_vlg_vec_tst is
end Circuit3_vlg_vec_tst;
