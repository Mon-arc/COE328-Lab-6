library verilog;
use verilog.vl_types.all;
entity Circuit2_vlg_vec_tst is
end Circuit2_vlg_vec_tst;
